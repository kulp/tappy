`default_nettype none
`timescale 10us/1us

module test(output clk, dat);

    initial
        $display("Starting test");

endmodule
